// emsys_alu : a simple ALU-like unit for the lab4 of the EmSys course 
//

module alu (
    input clk,
    input rst,

    // Inputs
	input logic [7:0] a,
	input logic [7:0] b,

	input logic [2:0] op,

    // Outputs
	output logic [7:0] q
);
// -------------------------------



endmodule

